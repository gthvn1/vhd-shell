conectix                 caml            `       `   �   �����c1��%B����{G�                                                                                                                                                                                                                                                                                                                                                                                                                                            cxsparse��������                 ���r                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������conectix                 caml            `       `   �   �����c1��%B����{G�                                                                                                                                                                                                                                                                                                                                                                                                                                            